//Created by Reetinder Kaur
//Modified by Nishant Mathur and Amanpreet Kaur
//Further Modified by Nishant Mathur
//Date 01 May 2017

//Changes from Lab 8 - 	1). DM & IM addr always available to mem_mod_mast irrespective of PL en. Now pipeline needs to be disabled and SW control enabled
//						2). All Dummies removed 
//						3). New signal SW ctrl added. refer mem_mod_mast for functionality
//						4). Data_mem_wea added as output from datapath
//						5). New signal PL done added to signal completion of instructions

//Changes from Lab 9 & Lab 10 -	1). Depth of Instruction memory has been increased from 512 locations to 4098 locations.

`timescale 1ns / 1ps

module datapath( clk,
				 rst,
				 pipeline_en,
				 sw_ctrl,
				 IorD,				// 1 for Data Memory
				 WorR,				// 1 for Read
				 
				 Addr_in,
				 Data_in,
				 IM_Addr_out,
				 DM_Addr_out,
				 IM_Data_out,
				 DM_Data_out,
				 
				 
				 EX_ALU_in1,
				 EX_ALU_in2,
				 EX_ALU_out,
				 EX_ALUop,
				
				 
				 RegWrite,
				 ALUSrc,
				 MemWrite,
				 MemtoReg,	
				 Jump,	
				 ble,	
				 imme,
				 ALUop,
				 PL_done,
				 FW_ld,
				 
				 Data_mem_dina,
				 Data_mem_addr,
				 Data_mem_wea, 
				 MEM_Dout, 
				 MEM_PL_done,
				 first_word
				);

//Inputs from Mem_mod_mast				
input clk;
input rst;
input pipeline_en;
input sw_ctrl;
input IorD;
input WorR;
input [8:0] Addr_in;
input [63:0] Data_in;
input [63:0] MEM_Dout;
input [7:0] first_word;
//input last_word;


//Control inputs from control

input RegWrite;
input ALUSrc;
input MemWrite;
input MemtoReg;	
input Jump;	
input ble;	
input imme; 
input [3:0] ALUop;
input PL_done;
input FW_ld;

//Output generated by ALU
input [63:0] EX_ALU_out;

//Data, address & control outputs to mem_mod_mast
output [8:0] IM_Addr_out;
output [8:0] DM_Addr_out;
output [31:0] IM_Data_out;
output [63:0] DM_Data_out;
output Data_mem_wea;
output [63:0] Data_mem_dina;
output [8:0] Data_mem_addr;
output MEM_PL_done;

//Inputs from EX to ALU
output [63:0] EX_ALU_in1, EX_ALU_in2;
output [3:0] EX_ALUop;



//reg [31:0] Dummy_data;
reg[8:0] IM_addra;
reg [31:0] IM_dina;
reg IM_wea;

//IF stage signals
wire [31:0] IF_Inst;
reg [8:0] IF_PC_out,IF_PC_out_next,IF_PC_out_after_thread_sel,IF_PC_out_next1,IF_PC_out_next2,IF_PC_out_next3,IF_PC_out_next4;
reg [1:0] thread_count,thread_count_next;

// ID stage signals
//reg ID_WRegEn, ID_WMemEn;
//reg [4:0] ID_Reg1, ID_Reg2;
//reg [4:0] ID_WReg1;
wire [63:0] ID_R1out, ID_R2out;
reg [63:0] ID_SGNEXT_val;
reg [8:0] ID_PC_out, Branch_Target,Branch_Offset;



// EX stage signals

reg EX_WRegEn, EX_WMemEn;
//reg [63:0] EX_R1out, EX_R2out;
//reg [55:0] EX_Dummy;
reg [4:0] EX_WReg1;
reg [63:0] EX_SGNEXT_val;
reg EX_ALUSrc, EX_MemtoReg;
reg PCSrc;
reg EX_ble, EX_Jump;
reg [8:0] EX_Branch_Target;
reg [3:0] EX_ALUop;
reg [63:0] EX_ALU_in1,EX_ALU_in2;
reg EX_PL_done;
reg EX_FW_ld;

// MEM stage signals
//reg Dummy_Addr;
reg [63:0] Data_mem_dina;
reg Data_mem_wea;
//reg [7:0] Data_mem_addra, Data_mem_addrb;
reg [7:0] Data_mem_addr;
reg MEM_WRegEn, MEM_WMemEn;
//reg [7:0] MEM_WAddr;
//reg [7:0] MEM_RAddr;
reg [63:0] MEM_ALU_out;
reg [63:0] MEM_Data;
reg [4:0] MEM_WReg1;
wire [63:0] MEM_Dout;
reg MEM_MemtoReg;
reg MEM_PL_done;
reg MEM_FW_ld;

// WB stage signals
reg WB_WRegEn;
//reg [63:0] WB_Dout;
reg [4:0] WB_WReg1;
reg [63:0] WB_ALUout;
reg [63:0] Reg_din,Reg_din_tmp;
reg WB_MemtoReg;
reg WB_FW_ld;

// Memory and Regfile instantiation
//data_mem data_mem(.clka(clk), .dina(Data_mem_dina),	.addra(Data_mem_addr), .wea(Data_mem_wea), .clkb(clk), .addrb(Data_mem_addr), .doutb(MEM_Dout)); -----removed for Lab 9 since intergration with convert FIFO carried out
inst_mem inst_mem(.clka(clk), .dina(IM_dina), .addra(IM_addra), .wea(IM_wea), .douta(IF_Inst));
regfile regfile(.clk(clk), .rst(rst), .r0addr(IF_Inst[19:15]), .r1addr(IF_Inst[24:20]), .waddr(WB_WReg1), .wdata(Reg_din), .wena(WB_WRegEn), .r0data(ID_R1out), .r1data(ID_R2out));

assign	IM_Addr_out = IM_addra;
assign	IM_Data_out = IF_Inst;
assign	DM_Addr_out = Data_mem_addr;
assign	DM_Data_out = MEM_Dout;


always @(posedge clk, posedge rst)
	begin
	
	if (rst == 1'b1)					//Reset entire pipeline
		begin
		IF_PC_out <= 9'h000;
		// IF_PC_out_after_thread_sel <= 'h0;
		// IF_PC_out_next1 <= 'h0;
		// IF_PC_out_next2 <= 'h7;
		// IF_PC_out_next3 <= 'hE;
		// IF_PC_out_next4 <= 'h15;
		thread_count <=2'b0;
//		ID_WRegEn <='h0;
//		ID_WMemEn <='h0;
//		ID_Reg1 <= 'h0;
//		ID_Reg2 <= 'h0;
//		ID_WReg1  <= 'h0;
		
		EX_WRegEn <= 'h0;
		EX_WMemEn <= 'h0;
//		EX_R1out <= 'h0;
//		EX_R2out <= 'h0;
		EX_WReg1 <= 'h0;
		EX_SGNEXT_val <= 'h0;
		EX_MemtoReg <= 'h0;
		EX_ALUSrc <= 'h0;
//		EX_PCSrc <= 'h0;
		EX_Branch_Target <= 'h0;
		EX_ALUop <= 'h0;
		EX_ble <= 'h0;
		EX_Jump <= 'h0;
		EX_PL_done <= 'h0;
		EX_FW_ld <= 'h0;
		
		MEM_WRegEn <= 'h0;
		MEM_WMemEn <= 'h0 ;
//		MEM_RAddr <= 'h0;
//		MEM_WAddr <= 'h0;
		MEM_ALU_out <= 'h0;
		MEM_Data <= 'h0 ;
		MEM_WReg1 <= 'h0 ;
		MEM_MemtoReg <= 'h0;
		MEM_PL_done <= 'h0;
		MEM_FW_ld <= 'h0;
		
//		WB_Dout <= 'h0 ;
		WB_WReg1 <= 'h0 ;
		WB_WRegEn <= 'h0 ;
		WB_ALUout <= 'h0;
		WB_MemtoReg <= 'h0;
		WB_FW_ld <= 'h0;
		
		end
	
	else if (pipeline_en == 1'b1 & IF_PC_out < 9'h120)
		begin
	
		// IF stage
		IF_PC_out <= IF_PC_out_next; 
		thread_count <= thread_count_next;
		
		
		
		// ID stage
//		ID_WRegEn <= RegWrite;							//RF write en
//		ID_WMemEn <= MemWrite;							//DM write en
//		ID_Reg1 <= IF_Inst[19:15];						//rs1 address
//		ID_Reg2 <= IF_Inst[24:20];						//rs2 address
//		ID_WReg1 <= IF_Inst[11:7];						//rd address
		ID_PC_out <= IF_PC_out;							//Carry PC value to ID stage
		
		
		// EX stage
		EX_WRegEn <= RegWrite;
		EX_WMemEn <= MemWrite;
//		EX_R1out <= ID_R1out;
//		EX_R2out <= ID_R2out;
		EX_WReg1 <= IF_Inst[11:7];
		EX_SGNEXT_val <= ID_SGNEXT_val;						//Carry sign extended immediate value or store address into EX
		EX_MemtoReg <= MemtoReg;							//Carry MemtoReg control signal to WB stage
		EX_ALUSrc <= ALUSrc;								//Carry ALUSrc to EX stage
//		EX_PCSrc <= PCSrc;									//Carry PCSrc to EX stage
		EX_Branch_Target <= Branch_Target;					//Carry Branch Target Address calculated to EX stage
		EX_ALUop <= ALUop;
		EX_Jump <= Jump;
		EX_ble <= ble;
		EX_PL_done <= PL_done;
		EX_FW_ld <= FW_ld;
		
		// MEM stage
		MEM_WRegEn <= EX_WRegEn ;
		MEM_WMemEn <= EX_WMemEn ;
		MEM_ALU_out <= EX_ALU_out;
//		MEM_RAddr <= EX_ALU_out[9:2];//EX_R1out[7:0] ;		//Addr calculted by ALU forwarded to D_MEM read port
//		EX_Dummy <= EX_ALU_out[63:10]//EX_R1out[63:8] ;		
//		MEM_WAddr <= EX_ALU_out[9:2];//EX_R1out[7:0] ;		//Addr calculted by ALU forwarded to D_MEM write port
		MEM_Data <= ID_R2out ;								//rs2 forwarded to MEM stage from before MUX
		MEM_WReg1 <= EX_WReg1 ;								//rd address
		MEM_MemtoReg <= EX_MemtoReg;						//Carry MemtoReg control signal to WB stage
		MEM_PL_done <= EX_PL_done;
		MEM_FW_ld <= EX_FW_ld;
		
		// WB stage
//		WB_Dout <= MEM_Dout;								//Give memory data out to WB stage
		WB_ALUout <= MEM_ALU_out;								//Give ALU calculated output to WB stage
		WB_WReg1 <= MEM_WReg1;								//rd address
		WB_WRegEn <= MEM_WRegEn;							//RF write en
		WB_MemtoReg <= MEM_MemtoReg;						//Carry MemtoReg control signal to WB stage
		WB_FW_ld <= MEM_FW_ld;
		
		
		end
		
	end

	always @(*)
	begin
	
	//IF stage controls and calculations

		
	//ID stage controls and calculations
	if (imme==1'b1)													//choose between ld/immediate values and store sign extended values 
		ID_SGNEXT_val = {{52{IF_Inst[31]}},IF_Inst[31:20]};
	else
		ID_SGNEXT_val = {{52{IF_Inst[31]}},IF_Inst[31:25],IF_Inst[11:7]};

	
	if (Jump)														//choose Branch_Offset based on jump/branch instruction
		Branch_Offset = IF_Inst[30:22];
	else
		Branch_Offset = {IF_Inst[30:25],IF_Inst[11:9]} ;
		
	Branch_Target = ID_PC_out + Branch_Offset;						//Calculate Branch Target
	
	//EX stage controls and calculations
//	EX_ALU_in1 = EX_R1out;		
	EX_ALU_in1 = ID_R1out;
	
	if (EX_ALUSrc)														//choose ALU src 2 from amongst rs2 and sign extended values 
		EX_ALU_in2 = EX_SGNEXT_val;										//Temprorary for testing
	else 
		EX_ALU_in2 = ID_R2out;
	
	if (EX_Jump | (EX_ble & ((ID_R1out == ID_R2out) | (ID_R2out < ID_R1out))))	//check for branch <= condition
		PCSrc = 'h1;
	else
		PCSrc = 'h0;
	
	if (MEM_PL_done || rst)
	begin
		IF_PC_out_after_thread_sel = 'h0;
		IF_PC_out_next1 = 'h0;
		IF_PC_out_next2 = 'h6;
		IF_PC_out_next3 = 'hD;
		IF_PC_out_next4 = 'h14;
		IF_PC_out_next = 'h0;
		thread_count_next = 'h0;
	end
	else if  (!(MEM_PL_done || rst) && pipeline_en)
	begin
	case(thread_count)
		'b00 : begin 
				IF_PC_out_next1=IF_PC_out;
				thread_count_next = 2'b01;
				IF_PC_out_after_thread_sel = IF_PC_out_next2 + 1;
//				IF_PC_out_after_thread_sel = IF_PC_out_next2;
				end
		'b01 : begin 
				IF_PC_out_next2=IF_PC_out;
				thread_count_next = 2'b10;
				IF_PC_out_after_thread_sel = IF_PC_out_next3 + 1;
//				IF_PC_out_after_thread_sel = IF_PC_out_next3;
				end
		'b10 : begin 
				IF_PC_out_next3=IF_PC_out;
				thread_count_next = 2'b11;
				IF_PC_out_after_thread_sel = IF_PC_out_next4 + 1;
//				IF_PC_out_after_thread_sel = IF_PC_out_next4;
				end
		'b11 : begin 
				IF_PC_out_next4=IF_PC_out;
				thread_count_next = 2'b00;
				IF_PC_out_after_thread_sel = IF_PC_out_next1 + 1;
//				IF_PC_out_after_thread_sel = IF_PC_out_next1;
				end
	endcase
	end
	else 
	begin
		IF_PC_out_next1 = IF_PC_out_next1;
		IF_PC_out_next2 = IF_PC_out_next2;
		IF_PC_out_next3 = IF_PC_out_next3;
		IF_PC_out_next4 = IF_PC_out_next4;
		thread_count_next = thread_count_next;
		IF_PC_out_after_thread_sel = IF_PC_out_after_thread_sel;

	end
	
	if (PCSrc)													//load PC value with branch target if branch condition is true, else increment PC
		IF_PC_out_next = EX_Branch_Target;
	else
		IF_PC_out_next = IF_PC_out_after_thread_sel;
		

		
	//MEM sstage memory initialization and address assignment
	//Set default vaues for IM & DM control, address and data pins
	IM_addra = IF_PC_out;  
	IM_wea = 1'b0;
	IM_dina = Data_in[31:0];
//	Dummy_data = Data_in[63:32];	
	
	Data_mem_dina = MEM_Data;
//	Data_mem_addrb = MEM_ALU_out[9:2];
//	Data_mem_addra = MEM_ALU_out[9:2];
	Data_mem_addr = MEM_ALU_out[9:2];
	Data_mem_wea = MEM_WMemEn;
	
		
	//Memory write and read access for user controlled arite and res operations from Mem_mod_mast
//	if (pipeline_en==1'b0)
//		begin
		if (!IorD)														//Write data to instruction and data memories based on ~I/D sel, pipeline en, write en and sw_ctrl
			begin
			if (!pipeline_en & sw_ctrl)
				begin
				IM_addra = Addr_in[8:0];
				if (!WorR)
					begin
//						IM_dina = Data_in[31:0];
						IM_wea = 'b1;
//						Dummy_data = Data_in[63:32]; 			
					end
				else	IM_wea = 1'b0;
				end
			end
		else
			begin
			if (!pipeline_en &  sw_ctrl)
				begin
				Data_mem_addr = Addr_in[7:0];
				if (!WorR)
					begin
//						Data_mem_addra = Addr_in[7:0];
						Data_mem_dina = Data_in;
						Data_mem_wea = 1'b1;
//						Dummy_Addr = Addr_in[8];
					end
				else	
					begin
//						Data_mem_addrb = Addr_in[7:0];
						Data_mem_wea = 1'b0;
//						Dummy_Addr = Addr_in[8];
					end
				end
			end
	
	//WB stage controls
	if (WB_FW_ld)
		Reg_din_tmp <= {first_word,2'b00};
	else
		Reg_din_tmp <= MEM_Dout;
	
	
	if (WB_MemtoReg)
			Reg_din	= WB_ALUout;					//Choose ALU calculated output or Memory Data output based (only for load instruction)
	else	
//			Reg_din	= WB_Dout;
			Reg_din	= Reg_din_tmp;
		
		
	end
endmodule












module datapath_tb;

reg clk, rst, pipeline_en, IorD, WorR;
reg [8:0] Addr_in;
reg [63:0] Data_in;
wire [8:0] IM_Addr_out, DM_Addr_out;
wire [63:0] DM_Data_out;
wire [31:0] IM_Data_out;
wire [63:0] EX_ALU_in1, EX_ALU_in2; 
reg [63:0] EX_ALU_out;
reg RegWrite, MemWrite, MemtoReg, Jump, ble, imme;
reg ALUSrc; 


// output clk, rst, pipeline_en, IorD, WorR; 
// output [8:0] Addr_in, 
// output [63:0] Data_in, 
// input [8:0] IM_Addr_out, 
// input [8:0] DM_Addr_out, 
// input [31:0] IM_Data_out, 
// input [63:0] DM_Data_out, 
// output [63:0] EX_ALU_in1, 
// output [63:0] EX_ALU_in2, 
// input [63:0] EX_ALU_out, 
// output RegWrite, ALUSrc, MemWrite,	 MemtoReg,	Jump, ble, imme;



datapath datapath(clk, rst, pipeline_en, IorD, WorR, Addr_in, Data_in, IM_Addr_out, DM_Addr_out, IM_Data_out, DM_Data_out, EX_ALU_in1, EX_ALU_in2, EX_ALU_out, RegWrite, ALUSrc, MemWrite,	 MemtoReg,	Jump, ble, imme);

initial
	begin
	rst=1;
	clk=0;
	pipeline_en=0;
	IorD=0;
	WorR=0;
	Addr_in=0;
	Data_in=0;
	RegWrite=0;
	ALUSrc=0;
	MemWrite=0;
	MemtoReg=0;
	Jump=0;
	ble=0;
	imme=0;
	
	forever #10 clk=~clk;	
	end

initial
	begin
	
	#9
	rst = 1'b0;		
	IorD=1'b1;
	WorR=1'b1;
	Addr_in=9'h000;
	
	#60
	RegWrite='h1;		//ld instruction
	ALUSrc = 'h1;
	imme = 'h1;
	
	
	
	
	#60
	Addr_in=9'h004;
	
	#60
	IorD=1'b0;
	WorR=1'b1;
	Addr_in=9'h000;
	
	#60
	Addr_in=9'h001;
	
	#60
	Addr_in=9'h002;
	
	#60
	pipeline_en=1'b1;
	
	#200
	pipeline_en=1'b0;
	IorD=1'b0;
	WorR=1'b0;
	Addr_in=9'h009;
	Data_in=64'hABCD12341234ABCD;
	
	#60
	IorD=1'b1;
	WorR=1'b0;
	Addr_in=9'h00C;
	Data_in=64'h12345678ABCDABCD;
	
	#60
	IorD=1'b0;
	WorR=1'b1;
	Addr_in=9'h009;
	
	#60
	IorD=1'b1;
	WorR=1'b1;
	Addr_in=9'h00C;
	
	end
				
endmodule 
